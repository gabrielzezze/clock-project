LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity divisor_generico is

generic (divisor : natural := 8);
    port(
      clk      :   in std_logic;
      saida_clk :   out std_logic;
		SW        :   in std_logic);

end entity;

-- O valor "n" do divisor, define a divisao por "2n".
-- Ou seja, n é metade do período da frequência de saída.

architecture div_inteiro of divisor_generico is

    signal tick : std_logic := '0';
    signal contador : integer range 0 to divisor+1 := 0;
	 signal divisor_inter : natural := divisor;

begin

	 divisor_inter <= divisor WHEN SW = '0' ELSE 250000;

    process(clk)
    begin
        if rising_edge(clk) then
            if contador = divisor_inter then
                contador <= 0;
                tick <= not tick;
            else
                contador <= contador + 1;
            end if;
        end if;
    end process;

saida_clk <= tick;

end architecture div_inteiro;
